`ifndef __MEMORY_SV
`define __MEMORY_SV

`ifdef VERILATOR
`include "include/common.sv"
`include "include/pipes.sv"
`include "pipeline/memory/read_data.sv"
`include "pipeline/memory/write_data.sv"
`else
`endif

module memory 
    import common::*;
    import pipes::*;(
    input logic clk,reset,
    input excute_data_t dataE,
    output memory_data_t dataM,
    output dbus_req_t  dreq,
	input  dbus_resp_t dresp,
    output logic stall_m,
    output forward_t forward_m
);
    
    msize_t msize;
    u1 mem_unsigned;
    word_t rslt,write_rslt,read_rslt;//result
    strobe_t strobe;
    always_comb begin
        unique case (dataE.ctl.op)
            LB,SB,LBU: msize=MSIZE1;
            LH,SH,LHU: msize=MSIZE2;
            LW,SW,LWU: msize=MSIZE4;
            LD,SD:     msize=MSIZE8;
            default: begin
                msize=MSIZE8;
            end 
        endcase
    end

    always_comb begin  
        unique case (dataE.ctl.op)
            LB,SB,LH,SH,LW,SW,LD,SD :mem_unsigned=0;
            LBU,LHU,LWU:mem_unsigned=1;
            default: begin
                mem_unsigned=0;
            end
        endcase
    end

    always_comb begin
        dreq='0;
        rslt=dataE.result;
        unique case(dataE.ctl.op)
            LB, LH, LW, LBU, LHU, LWU, LD: begin
                dreq.valid=dataE.valid;
                dreq.addr=dataE.result;
                dreq.size=msize;
                
                rslt=read_rslt;      
            end
            SB, SH, SW, SD: begin
                dreq.valid=dataE.valid;
                dreq.addr=dataE.result;
                dreq.size=msize;
                dreq.strobe=strobe;
                dreq.data=write_rslt;     
            end
            default: begin
                
            end
        endcase
    end
    read_data read_data(
        ._rd(dresp.data),.rd(read_rslt),
        .addr(dataE.result[2:0]),
        .msize,.mem_unsigned
    );
    write_data write_data(
        ._wd(dataE.rd2),.wd(write_rslt),
        .addr(dataE.result[2:0]),
        .msize,.strobe
    );

    logic bubble;

    always_comb begin
    unique case(dataE.ctl.op)
        LB, LH, LW, LBU, LHU, LWU, LD,
        SB, SH, SW, SD:
            bubble=~dresp.data_ok; 
        default: 
            bubble = 0;
        endcase
    end

    assign stall_m=bubble&(dataE.valid);
    //only needs to be paused when a valid instr is processed
    //and the memory op is not completed

    assign forward_m.dst=(dataE.ctl.regwrite & dataE.valid)?dataE.dst:0;
    assign forward_m.data=rslt;
    assign forward_m.ismem=1;

    always_ff @(posedge clk) begin
        if (reset) begin
            dataM.valid <= 0;
        end else begin
            if (stall_m) dataM.valid<=0;
            else begin
                dataM.pc <= dataE.pc;
                dataM.valid <= dataE.valid;
                dataM.raw_instr <= dataE.raw_instr;
                dataM.result <= rslt;
                dataM.ctl <= dataE.ctl;
                dataM.dst <= dataE.dst; 
                dataM.addr <= dataE.result;
            end
        end
    end


endmodule
`endif